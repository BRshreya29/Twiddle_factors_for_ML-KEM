`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 24.01.2025 23:50:07
// Design Name: 
// Module Name: twiddlefactor_storage_unit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module store_phi_values (
    input [7:0] p,   // 8-bit input for p (0 to 255)
    output reg [11:0] phi // 12-bit output for phi values
);
    always @(*) begin
        case (p)
        8'd0   : phi = 12'd1;
8'd1   : phi = 12'd2688;
8'd2   : phi = 12'd1414;
8'd3   : phi = 12'd2443;
8'd4   : phi = 12'd1996;
8'd5   : phi = 12'd2229;
8'd6   : phi = 12'd2681;
8'd7   : phi = 12'd2572;
8'd8   : phi = 12'd2532;
8'd9   : phi = 12'd1540;
8'd10  : phi = 12'd1573;
8'd11  : phi = 12'd394;
8'd12  : phi = 12'd450;
8'd13  : phi = 12'd1173;
8'd14  : phi = 12'd461;
8'd15  : phi = 12'd780;
8'd16  : phi = 12'd2699;
8'd17  : phi = 12'd1021;
8'd18  : phi = 12'd1352;
8'd19  : phi = 12'd2237;
8'd20  : phi = 12'd882;
8'd21  : phi = 12'd568;
8'd22  : phi = 12'd2102;
8'd23  : phi = 12'd863;
8'd24  : phi = 12'd2760;
8'd25  : phi = 12'd1868;
8'd26  : phi = 12'd1052;
8'd27  : phi = 12'd1455;
8'd28  : phi = 12'd2794;
8'd29  : phi = 12'd48;
8'd30  : phi = 12'd2522;
8'd31  : phi = 12'd1292;
8'd32  : phi = 12'd749;
8'd33  : phi = 12'd2596;
8'd34  : phi = 12'd464;
8'd35  : phi = 12'd2186;
8'd36  : phi = 12'd283;
8'd37  : phi = 12'd1692;
8'd38  : phi = 12'd682;
8'd39  : phi = 12'd2266;
8'd40  : phi = 12'd2267;
8'd41  : phi = 12'd1626;
8'd42  : phi = 12'd3040;
8'd43  : phi = 12'd2154;
8'd44  : phi = 12'd821;
8'd45  : phi = 12'd3050;
8'd46  : phi = 12'd2402;
8'd47  : phi = 12'd1645;
8'd48  : phi = 12'd848;
8'd49  : phi = 12'd2388;
8'd50  : phi = 12'd632;
8'd51  : phi = 12'd1026;
8'd52  : phi = 12'd1476;
8'd53  : phi = 12'd2649;
8'd54  : phi = 12'd3110;
8'd55  : phi = 12'd561;
8'd56  : phi = 12'd3260;
8'd57  : phi = 12'd952;
8'd58  : phi = 12'd2304;
8'd59  : phi = 12'd1212;
8'd60  : phi = 12'd2094;
8'd61  : phi = 12'd2662;
8'd62  : phi = 12'd1435;
8'd63  : phi = 12'd2298;
8'd64  : phi = 12'd1729;
8'd65  : phi = 12'd268;
8'd66  : phi = 12'd1320;
8'd67  : phi = 12'd2775;
8'd68  : phi = 12'd2240;
8'd69  : phi = 12'd2288;
8'd70  : phi = 12'd1481;
8'd71  : phi = 12'd2773;
8'd72  : phi = 12'd193;
8'd73  : phi = 12'd2789;
8'd74  : phi = 12'd3253;
8'd75  : phi = 12'd2110;
8'd76  : phi = 12'd2393;
8'd77  : phi = 12'd756;
8'd78  : phi = 12'd1438;
8'd79  : phi = 12'd375;
8'd80  : phi = 12'd2642;
8'd81  : phi = 12'd939;
8'd82  : phi = 12'd650;
8'd83  : phi = 12'd2804;
8'd84  : phi = 12'd296;
8'd85  : phi = 12'd17;
8'd86  : phi = 12'd2419;
8'd87  : phi = 12'd735;
8'd88  : phi = 12'd1583;
8'd89  : phi = 12'd642;
8'd90  : phi = 12'd1274;
8'd91  : phi = 12'd2300;
8'd92  : phi = 12'd447;
8'd93  : phi = 12'd3096;
8'd94  : phi = 12'd2877;
8'd95  : phi = 12'd109;
8'd96  : phi = 12'd40;
8'd97  : phi = 12'd992;
8'd98  : phi = 12'd3296;
8'd99  : phi = 12'd1179;
8'd100 : phi = 12'd3273;
8'd101 : phi = 12'd2606;
8'd102 : phi = 12'd712;
8'd103 : phi = 12'd3010;
8'd104 : phi = 12'd1410;
8'd105 : phi = 12'd1678;
8'd106 : phi = 12'd2998;
8'd107 : phi = 12'd2444;
8'd108 : phi = 12'd1355;
8'd109 : phi = 12'd314;
8'd110 : phi = 12'd1795;
8'd111 : phi = 12'd1239;
8'd112 : phi = 12'd1432;
8'd113 : phi = 12'd892;
8'd114 : phi = 12'd816;
8'd115 : phi = 12'd2926;
8'd116 : phi = 12'd1990;
8'd117 : phi = 12'd2746;
8'd118 : phi = 12'd855;
8'd119 : phi = 12'd1230;
8'd120 : phi = 12'd543;
8'd121 : phi = 12'd1482;
8'd122 : phi = 12'd2132;
8'd123 : phi = 12'd1607;
8'd124 : phi = 12'd1903;
8'd125 : phi = 12'd1920;
8'd126 : phi = 12'd1010;
8'd127 : phi = 12'd1745;

            
                      8'd128 : phi = 12'd660;
8'd129 : phi = 12'd1881;
8'd130 : phi = 12'd1226;
8'd131 : phi = 12'd3022;
8'd132 : phi = 12'd2404;
8'd133 : phi = 12'd1129;
8'd134 : phi = 12'd1882;
8'd135 : phi = 12'd2938;
8'd136 : phi = 12'd1305;
8'd137 : phi = 12'd2603;
8'd138 : phi = 12'd2764;
8'd139 : phi = 12'd2657;
8'd140 : phi = 12'd120;
8'd141 : phi = 12'd1665;
8'd142 : phi = 12'd1277;
8'd143 : phi = 12'd2246;
8'd144 : phi = 12'd1396;
8'd145 : phi = 12'd2584;
8'd146 : phi = 12'd2737;
8'd147 : phi = 12'd2148;
8'd148 : phi = 12'd2885;
8'd149 : phi = 12'd1557;
8'd150 : phi = 12'd1039;
8'd151 : phi = 12'd222;
8'd152 : phi = 12'd1484;
8'd153 : phi = 12'd1425;
8'd154 : phi = 12'd3313;
8'd155 : phi = 12'd1984;
8'd156 : phi = 12'd3028;
8'd157 : phi = 12'd305;
8'd158 : phi = 12'd1764;
8'd159 : phi = 12'd2791;
8'd160 : phi = 12'd826;
8'd161 : phi = 12'd3087;
8'd162 : phi = 12'd1310;
8'd163 : phi = 12'd1342;
8'd164 : phi = 12'd1968;
8'd165 : phi = 12'd2438;
8'd166 : phi = 12'd210;
8'd167 : phi = 12'd2449;
8'd168 : phi = 12'd231;
8'd169 : phi = 12'd2089;
8'd170 : phi = 12'd2116;
8'd171 : phi = 12'd2592;
8'd172 : phi = 12'd3168;
8'd173 : phi = 12'd2620;
8'd174 : phi = 12'd2447;
8'd175 : phi = 12'd1727;
8'd176 : phi = 12'd2579;
8'd177 : phi = 12'd3163;
8'd178 : phi = 12'd3223;
8'd179 : phi = 12'd3186;
8'd180 : phi = 12'd2242;
8'd181 : phi = 12'd695;
8'd182 : phi = 12'd344;
8'd183 : phi = 12'd3245;
8'd184 : phi = 12'd3122;
8'd185 : phi = 12'd877;
8'd186 : phi = 12'd186;
8'd187 : phi = 12'd1852;
8'd188 : phi = 12'd2083;
8'd189 : phi = 12'd277;
8'd190 : phi = 12'd1752;
8'd191 : phi = 12'd1377;
8'd192 : phi = 12'd1333;
8'd193 : phi = 12'd2502;
8'd194 : phi = 12'd312;
8'd195 : phi = 12'd1154;
8'd196 : phi = 12'd2881;
8'd197 : phi = 12'd264;
8'd198 : phi = 12'd135;
8'd199 : phi = 12'd1020;
8'd200 : phi = 12'd2490;
8'd201 : phi = 12'd3106;
8'd202 : phi = 12'd1366;
8'd203 : phi = 12'd1981;
8'd204 : phi = 12'd1887;
8'd205 : phi = 12'd1370;
8'd206 : phi = 12'd2158;
8'd207 : phi = 12'd287;
8'd208 : phi = 12'd1576;
8'd209 : phi = 12'd2292;
8'd210 : phi = 12'd288;
8'd211 : phi = 12'd2695;
8'd212 : phi = 12'd3000;
8'd213 : phi = 12'd1486;
8'd214 : phi = 12'd2414;
8'd215 : phi = 12'd1124;
8'd216 : phi = 12'd2328;
8'd217 : phi = 12'd3052;
8'd218 : phi = 12'd900;
8'd219 : phi = 12'd1718;
8'd220 : phi = 12'd1523;
8'd221 : phi = 12'd466;
8'd222 : phi = 12'd2675;
8'd223 : phi = 12'd1050;
8'd224 : phi = 12'd733;
8'd225 : phi = 12'd1726;
8'd226 : phi = 12'd3243;
8'd227 : phi = 12'd2078;
8'd228 : phi = 12'd1118;
8'd229 : phi = 12'd2111;
8'd230 : phi = 12'd2982;
8'd231 : phi = 12'd2901;
8'd232 : phi = 12'd1198;
8'd233 : phi = 12'd1257;
8'd234 : phi = 12'd1371;
8'd235 : phi = 12'd2063;
8'd236 : phi = 12'd2685;
8'd237 : phi = 12'd1358;
8'd238 : phi = 12'd1126;
8'd239 : phi = 12'd1560;
8'd240 : phi = 12'd3183;
8'd241 : phi = 12'd3257;
8'd242 : phi = 12'd2876;
8'd243 : phi = 12'd2173;
8'd244 : phi = 12'd1041;
8'd245 : phi = 12'd1042;
8'd246 : phi = 12'd2374;
8'd247 : phi = 12'd1291;
8'd248 : phi = 12'd3234;
8'd249 : phi = 12'd153;
8'd250 : phi = 12'd3254;
8'd251 : phi = 12'd947;
8'd252 : phi = 12'd2371;
8'd253 : phi = 12'd2717;
8'd254 : phi = 12'd1461;
8'd255 : phi = 12'd0;


        endcase
    end
endmodule